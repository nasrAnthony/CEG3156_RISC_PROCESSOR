library ieee;
use ieee.std_logic_1164.all;

entity decode3t8 is 
	port 
		(
		);
end entity;


architecture struct of decode3t8 is 
signal int_inp : std_logic_vector(7 downto 0);
