instrMemoryREG_inst : instrMemoryREG PORT MAP (
		address	 => address_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
